
package vsc_tr;

endpackage
